interface Intf();
	`debug
endinterface
