interface Intf();
endinterface
