`ifndef envPkg__sv
`define envPkg__sv

package envPkg;
	`include "uvm_macros.svh"
	import uvm_pkg::*;
	import rhudbg::*;

	`include "baseTest.svh"

endpackage
`endif
